-------------------------------------------------------------------------------
-- Project     : audio_top
-- Description : Constants and LUT for tone generation with DDS
--
--
-------------------------------------------------------------------------------
--
-- Change History
-- Date     |Name      |Modification
------------|----------|-------------------------------------------------------
-- 12.04.13 | dqtm     | file created for DTP2 Milestone-3 in FS13
-- 02.04.14 | dqtm     | updated for DTP2 in FS14, cause using new parameters
-- 27.04.18 | dqtm     | updated for EA999 in FS18, check naming compatibility with filter_pkg
-------------------------------------------------------------------------------

-------------------------------------------------------------------------------
-- Package  Declaration
-------------------------------------------------------------------------------
-- Include in Design of Block dds.vhd and tone_decoder.vhd :
--   use work.tone_gen_pkg.all;
-------------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package DSVF_pkg is


    -------------------------------------------------------------------------------
	-- CONSTANT DECLARATION FOR SEVERAL BLOCKS
	-------------------------------------------------------------------------------


	constant N_DATA_HALF_RESOL		: natural := 8;
	constant N_DATA_RESOL			: natural := 16;			-- data Bus width (MSB determina sinal)
	constant N_DATA_DOUBLE_RESOL 	: natural := 32;
	constant N_DATA_RESOL_WS 		: natural := 24; 
	constant N_MIDI_DATA 			: natural := 7;			-- number of data bits in MIDI mensage
	constant L_MIDI 					: natural := 2**N_MIDI_DATA; 
	-------------------------------------------------------------------------------
	-- TYPE DECLARATION FOR DDS
	-------------------------------------------------------------------------------
    subtype t_filter_range is integer range 0 to (65536);  -- range : [0; (2^16)]

	type filter_lut_rom is array (0 to L_MIDI-1) of t_filter_range;

	constant LUT_freq : filter_lut_rom := (
	1085,1115,1146,1177,1210,1243,1277,1313,1349,1386,1424,1463,1504,
	1545,1588,1632,1677,1723,1770,1819,1869,1921,1974,2028,2084,2141,
	2200,2261,2323,2387,2453,2521,2590,2661,2735,2810,2888,2967,3049,
	3133,3219,3308,3399,3493,3589,3688,3789,3894,4001,4111,4224,4340,
	4460,4583,4709,4838,4971,5108,5249,5393,5541,5694,5850,6011,6176,
	6346,6521,6700,6884,7073,7267,7467,7671,7882,8098,8320,8548,8783,
	9023,9270,9524,9785,10052,10327,10609,10899,11197,11502,11816,12138,
	12469,12808,13156,13514,13881,14257,14644,15040,15447,15865,16293,
	16732,17183,17645,18119,18605,19103,19613,20137,20673,21222,21785,
	22362,22952,23556,24175,24808,25456,26118,26796,27489,28197,28920,
	29659,30413,31182,31967,32768 );
	
	constant LUT_resson : filter_lut_rom := (
	48467,46429,44476,42606,40814,39097,37453,35877,34368,32923,31538,
	30212,28941,27724,26558,25441,24371,23346,22364,21423,20522,19659,
	18832,18040,17281,16554,15858,15191,14552,13940,13354,12792,12254,
	11739,11245,10772,10319,9885,9469,9071,8689,8324,7974,7639,7317,
	7009,6715,6432,6162,5903,5654,5416,5189,4970,4761,4561,4369,4186,
	4009,3841,3679,3525,3376,3234,3098,2968,2843,2724,2609,2499,2394,
	2293,2197,2105,2016,1931,1850,1772,1698,1626,1558,1492,1430,1369,
	1312,1257,1204,1153,1105,1058,1014,971,930,891,854,818,783,750,719,
	689,660,632,605,580,555,532,510,488,468,448,429,411,394,377,361,346,
	332,318,304,292,279,268,256,246,235,225,216,207 );
	
	-- 32 equivale ao valor 1 em Q3.5
    constant LUT_gain : filter_lut_rom := (
    1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,
    27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,
    50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,
    73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,
    96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,
    114,115,116,117,118,119,120,121,122,123,124,125,126,127,128 );
	
	constant LUT_waveshaping : filter_lut_rom := (
	4915,4966,5017,5067,5116,5166,5215,5264,5312,5360,5408,5456,5502,5549,
	5595,5641,5686,5731,5775,5819,5862,5905,5947,5989,6031,6071,6112,6152,
	6191,6230,6268,6306,6343,6380,6416,6452,6487,6522,6556,6589,6622,6655,
	6687,6719,6749,6780,6810,6839,6868,6897,6925,6952,6979,7006,7032,7057,
	7082,7107,7131,7154,7178,7200,7223,7245,7266,7287,7308,7328,7348,7367,
	7386,7405,7423,7441,7458,7475,7492,7508,7524,7540,7555,7570,7585,7599,
	7613,7627,7641,7654,7667,7679,7692,7704,7715,7727,7738,7749,7760,7770,
	7780,7790,7800,7810,7819,7828,7837,7846,7854,7862,7870,7878,7886,7894,
	7901,7908,7915,7922,7929,7935,7941,7948,7954,7960,7965,7971,7976,7982,
	7987,7992 );
	-------------------------------------------------------------------------------		
end package;
